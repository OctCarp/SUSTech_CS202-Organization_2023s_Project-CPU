`ifndef _VGA_HEAD
`define _VGA_HEAD

`timescale 1ps / 1ps

parameter _v0 = 6'b00_0000;
parameter _v1 = 6'b00_0001;
parameter _v2 = 6'b00_0010;
parameter _v3 = 6'b00_0011;
parameter _v4 = 6'b00_0100;
parameter _v5 = 6'b00_0101;
parameter _v6 = 6'b00_0110;
parameter _v7 = 6'b00_0111;
parameter _v8 = 6'b00_1000;
parameter _v9 = 6'b00_1001;


parameter _vA = 6'b00_1010;
parameter _vB = 6'b00_1011;
parameter _vC = 6'b00_1100;
parameter _vD = 6'b00_1101;
parameter _vE = 6'b00_1110;
parameter _vF = 6'b00_1111;
parameter _vG = 6'b01_0000;
parameter _vH = 6'b01_0001;
parameter _vI = 6'b01_0010;
parameter _vJ = 6'b01_0011;
parameter _vK = 6'b01_0100;
parameter _vL = 6'b01_0101;
parameter _vM = 6'b01_0110;
parameter _vN = 6'b01_0111;
parameter _vO = 6'b01_1000;
parameter _vP = 6'b01_1001;
parameter _vQ = 6'b01_1010;
parameter _vR = 6'b01_1011;
parameter _vS = 6'b01_1100;
parameter _vT = 6'b01_1101;
parameter _vU = 6'b01_1110;
parameter _vV = 6'b01_1111;
parameter _vW = 6'b10_0000;
parameter _vX = 6'b10_0001;
parameter _vY = 6'b10_0010;
parameter _vZ = 6'b10_0011;

parameter _SLASH = 6'b10_0100;
parameter _SPACE = 6'b11_1110;
parameter _COLON = 6'b11_1111;

`endif
